-------------------------------------------------------------------------
-- Group 9
-- Project Part A 
-- Lab Date: 09/28/11 +10/5/2011
-------------------------------------------------------------------------

-- tb_ALU32.vhd
-------------------------------------------------------------------------
-- DESCRIPTION:  This is a testbench to test our 32 bit ALU 
--
-------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;
use WORK.mips_package.all;

entity tb_ALU32 is

end tb_ALU32;

architecture behavioral of tb_ALU32 is


Component ALU32 is
  port(i_A       : in std_logic_vector(31 downto 0);
       i_B       : in std_logic_vector(31 downto 0);
       i_Opcode  : in std_logic_vector(2 downto 0);
       o_F       : out std_logic_vector(31 downto 0);
       o_CryOut  : out std_logic;
       o_Overflow: out std_logic;
       o_Zero    : out std_logic);

end Component;



signal s_A, s_B, s_F                        : std_logic_vector(31 downto 0);
signal s_Opcode                             : std_logic_vector(2 downto 0);
signal s_Zero, s_Overflow, s_CryOut         : std_logic;

begin
  testme: ALU32 

  port map(i_A => s_A,
           i_B => s_B,
           i_Opcode => s_Opcode,
           o_F => s_F,
           o_CryOut => s_CryOut,
           o_Overflow => s_Overflow,
           o_Zero => s_Zero);
  	        
  
process
begin


-------------------------------------------------------------------------
-- And test !!!!!
--  
--
-- This will test our and function of our 32 bit ALU
--
--
--And Test
-------------------------------------------------------------------------

-------------------------------------------------------------------------
-- 0 and 0
-- Expected value F= x000000000, CryOut= 0, Zero= 1,  overFlow =0
-------------------------------------------------------------------------

    s_A <= x"00000000";
    s_B <= x"00000000";
    s_Opcode <= "000";
    wait for 100 ns;

-------------------------------------------------------------------------
-- 1 and 1
-- Expected value F= x000000001, CryOut= 0, Zero= 0,  overFlow =0
-------------------------------------------------------------------------

    s_A <= x"00000001";
    s_B <= x"00000001";
    s_Opcode <= "000";
    wait for 100 ns;

-------------------------------------------------------------------------
-- 00000000 and FFFFFFFF
-- Expected value F= x000000000, CryOut= 0, Zero= 1,  overFlow =0
-------------------------------------------------------------------------

    s_A <= x"00000000";
    s_B <= x"FFFFFFFF";
    s_Opcode <= "000";
    wait for 100 ns;

-------------------------------------------------------------------------
-- FFFFFFFF and FFFFFFFF
-- Expected value F= xFFFFFFFF, CryOut= 0, Zero= 0,  overFlow =0
-------------------------------------------------------------------------

    s_A <= x"FFFFFFFF";
    s_B <= x"FFFFFFFF";
    s_Opcode <= "000";
    wait for 100 ns;




-------------------------------------------------------------------------
-- End of And test !!!!!
--  
--
-- 
--
--
--End of And Test
-------------------------------------------------------------------------



-------------------------------------------------------------------------
-- Or test !!!!!
--  
--
-- This will test our or function of our 32 bit ALU
--
--
--OR Test
-------------------------------------------------------------------------

-------------------------------------------------------------------------
-- 0 or 0
-- Expected value F= x000000000, CryOut= 0, Zero= 1,  overFlow =0
-------------------------------------------------------------------------

    s_A <= x"00000000";
    s_B <= x"00000000";
    s_Opcode <= "001";
    wait for 100 ns;

-------------------------------------------------------------------------
-- 0 or 1
-- Expected value F= x00000001, CryOut= 0, Zero= 0,  overFlow =0
-------------------------------------------------------------------------

    s_A <= x"00000000";
    s_B <= x"00000001";
    s_Opcode <= "001";
    wait for 100 ns;

-------------------------------------------------------------------------
-- 00000000 or FFFFFFFF
-- Expected value F= xFFFFFFFF, CryOut= 0, Zero= 0,  overFlow =0
-------------------------------------------------------------------------

    s_A <= x"00000000";
    s_B <= x"FFFFFFFF";
    s_Opcode <= "001";
    wait for 100 ns;

-------------------------------------------------------------------------
-- FFFFFFFF or 00000000  
-- Expected value F= xFFFFFFFF, CryOut= 0, Zero= 0,  overFlow =0
-------------------------------------------------------------------------

    s_A <= x"FFFFFFFF";
    s_B <= x"00000000";
    s_Opcode <= "001";
    wait for 100 ns;


-------------------------------------------------------------------------
-- FFFFFFFF or FFFFFFFF 
-- Expected value F= xFFFFFFFF, CryOut= 0, Zero= 0,  overFlow =0
-------------------------------------------------------------------------

    s_A <= x"FFFFFFFF";
    s_B <= x"FFFFFFFF";
    s_Opcode <= "001";
    wait for 100 ns;

-------------------------------------------------------------------------
-- End   Or test !!!!!
--  
--
-- 
--
--
-- End OR Test !!!!!!!!!
-------------------------------------------------------------------------

-------------------------------------------------------------------------
-- xor test !!!!!
--  
--
-- This will test our xor function of our 32 bit ALU
--
--
-- xor Test
-------------------------------------------------------------------------

-------------------------------------------------------------------------
-- 00000000 xor 00000000 
-- Expected value F= x00000000, CryOut= 0, Zero= 1,  overFlow =0
-------------------------------------------------------------------------

    s_A <= x"00000000";
    s_B <= x"00000000";
    s_Opcode <= "010";
    wait for 100 ns;

-------------------------------------------------------------------------
-- FFFFFFFF xor 00000000 
-- Expected value F= xFFFFFFFF, CryOut= 0, Zero= 0,  overFlow =0
-------------------------------------------------------------------------

    s_A <= x"FFFFFFFF";
    s_B <= x"00000000";
    s_Opcode <= "010";
    wait for 100 ns;
    
-------------------------------------------------------------------------
-- 00000000 xor FFFFFFFF 
-- Expected value F= xFFFFFFFF, CryOut= 0, Zero= 0,  overFlow =0
-------------------------------------------------------------------------

    s_A <= x"00000000";
    s_B <= x"FFFFFFFF";
    s_Opcode <= "010";
    wait for 100 ns;
    
-------------------------------------------------------------------------
-- FFFFFFFF xor FFFFFFFF 
-- Expected value F= x00000000, CryOut= 0, Zero= 1,  overFlow =0
-------------------------------------------------------------------------

    s_A <= x"FFFFFFFF";
    s_B <= x"FFFFFFFF";
    s_Opcode <= "010";
    wait for 100 ns;   

-------------------------------------------------------------------------
-- End   xOr test !!!!!
--  
--
-- 
--
--
-- End XOR Test !!!!!!!!!
-------------------------------------------------------------------------

-------------------------------------------------------------------------
-- nand test !!!!!
--  
--
-- This will test our nand function of our 32 bit ALU
--
--
--nand Test
-------------------------------------------------------------------------

-------------------------------------------------------------------------
-- 00000000 nand 00000000 
-- Expected value F= xFFFFFFFF, CryOut= 0, Zero= 0,  overFlow =0
-------------------------------------------------------------------------

    s_A <= x"00000000";
    s_B <= x"00000000";
    s_Opcode <= "011";
    wait for 100 ns;
    
-------------------------------------------------------------------------
-- FFFFFFFF nand 00000000 
-- Expected value F= xFFFFFFFF, CryOut= 0, Zero= 0,  overFlow =0
-------------------------------------------------------------------------

    s_A <= x"FFFFFFFF";
    s_B <= x"00000000";
    s_Opcode <= "011";
    wait for 100 ns;
 
-------------------------------------------------------------------------
-- 00000000 nand FFFFFFFF
-- Expected value F= xFFFFFFFF, CryOut= 0, Zero= 0,  overFlow =0
-------------------------------------------------------------------------

    s_A <= x"00000000";
    s_B <= x"FFFFFFFF";
    s_Opcode <= "011";
    wait for 100 ns;  
    
-------------------------------------------------------------------------
-- FFFFFFFF nand FFFFFFFF 
-- Expected value F= x00000000, CryOut= 0, Zero= 1,  overFlow =0
-------------------------------------------------------------------------

    s_A <= x"FFFFFFFF";
    s_B <= x"FFFFFFFF";
    s_Opcode <= "011";
    wait for 100 ns;
    

-------------------------------------------------------------------------
-- End  nand test !!!!!
--  
--
-- 
--
--
-- End NAND Test !!!!!!!!!
-------------------------------------------------------------------------

-------------------------------------------------------------------------
-- nor test !!!!!
--  
--
-- This will test our nor function of our 32 bit ALU
--
--
--nor Test
-------------------------------------------------------------------------

-------------------------------------------------------------------------
-- 00000000 nor 00000000 
-- Expected value F= xFFFFFFFF, CryOut= 0, Zero= 0,  overFlow =0
-------------------------------------------------------------------------

    s_A <= x"00000000";
    s_B <= x"00000000";
    s_Opcode <= "100";
    wait for 100 ns;

-------------------------------------------------------------------------
-- FFFFFFFF nor 00000000 
-- Expected value F= x00000000, CryOut= 0, Zero= 1,  overFlow =0
-------------------------------------------------------------------------

    s_A <= x"FFFFFFFF";
    s_B <= x"00000000";
    s_Opcode <= "100";
    wait for 100 ns;
    
-------------------------------------------------------------------------
-- 00000000 nor FFFFFFFF 
-- Expected value F= x00000000, CryOut= 0, Zero= 1,  overFlow =0
-------------------------------------------------------------------------

    s_A <= x"00000000";
    s_B <= x"FFFFFFFF";
    s_Opcode <= "100";
    wait for 100 ns;
    
-------------------------------------------------------------------------
-- FFFFFFFF nor FFFFFFFF 
-- Expected value F= x00000000, CryOut= 0, Zero= 1,  overFlow =0
-------------------------------------------------------------------------

    s_A <= x"FFFFFFFF";
    s_B <= x"FFFFFFFF";
    s_Opcode <= "100";
    wait for 100 ns;   
  
-------------------------------------------------------------------------
-- End  nor test !!!!!
--  
--
-- 
--
--
-- End NOR Test !!!!!!!!!
-------------------------------------------------------------------------
 
  
-------------------------------------------------------------------------
-- Add test !!!!!
--  
--
-- This will test our add function of our 32 bit ALU
--
--
--Add Test
-------------------------------------------------------------------------

-------------------------------------------------------------------------
-- 0 + 0
-- Expected value F= 0, CryOut= 0, Zero= 1,  overFlow =0
-------------------------------------------------------------------------
    s_A <= x"00000000";
    s_B <= x"00000000";
    s_Opcode <= "101";
    wait for 100 ns;
 
-------------------------------------------------------------------------
-- 0 + 1
-- Expected value F= 1, CryOut= 0, Zero= 0,  overFlow =0
-------------------------------------------------------------------------
    s_A <= x"00000000";
    s_B <= x"00000001";
    s_Opcode <= "101";
    wait for 100 ns; 
    
-------------------------------------------------------------------------
--  0 + -5
-- Expected value F= -5, CryOut= 0, Zero= 0,  overFlow =0
-------------------------------------------------------------------------
    s_A <= x"00000000";
    s_B <= x"FFFFFFFB";
    s_Opcode <= "101";
    wait for 100 ns;   

    
-------------------------------------------------------------------------
--  6 + -5
-- Expected value F= 1, CryOut= 1, Zero= 0,  overFlow =0
-------------------------------------------------------------------------
    s_A <= x"00000006";
    s_B <= x"FFFFFFFB";
    s_Opcode <= "101";
    wait for 100 ns;   
    
-------------------------------------------------------------------------
--  1 + 2147483647
-- Expected value F= 80000000, CryOut= 1, Zero= 0,  overFlow =1
-------------------------------------------------------------------------
    s_A <= x"7FFFFFFF";
    s_B <= x"00000001";
    s_Opcode <= "101";
    wait for 100 ns;   
  
-------------------------------------------------------------------------
-- End of Add test !!!!!
--  
--
-- 
--
--
--End of Add Test !!!!!!
-------------------------------------------------------------------------   

-------------------------------------------------------------------------
-- SLT test !!!!!
--  
--
-- This will test our SLT function of our 32 bit ALU
--
--
--SLT Test
-------------------------------------------------------------------------

-------------------------------------------------------------------------
-- 0 < 0
-- Expected value F= x00000000, CryOut= 0, Zero= 1,  overFlow =0
-------------------------------------------------------------------------
    s_A <= x"00000000";
    s_B <= x"00000000";
    s_Opcode <= "110";
    wait for 100 ns;

-------------------------------------------------------------------------
-- 1 < 0
-- Expected value F= x00000000, CryOut= 0, Zero= 1,  overFlow =0
-------------------------------------------------------------------------
    s_A <= x"00000001";
    s_B <= x"00000000";
    s_Opcode <= "110";
    wait for 100 ns;    
    
-------------------------------------------------------------------------
-- 1 < 2
-- Expected value F= x00000001, CryOut= 0, Zero= 0,  overFlow =0
-------------------------------------------------------------------------
    s_A <= x"00000001";
    s_B <= x"00000002";
    s_Opcode <= "110";
    wait for 100 ns; 
    
    
-------------------------------------------------------------------------
-- FFFFFFFF < 0
-- Expected value F= x00000001, CryOut= 0, Zero= 0,  overFlow =0
-------------------------------------------------------------------------
    s_A <= x"FFFFFFFF";
    s_B <= x"00000000";
    s_Opcode <= "110";
    wait for 100 ns;
    
-------------------------------------------------------------------------
-- 00000000 < FFFFFFFF
-- Expected value F= x00000000, CryOut= 0, Zero= 1,  overFlow =0
-------------------------------------------------------------------------
    s_A <= x"FFFFFFFF";
    s_B <= x"00000000";
    s_Opcode <= "110";
    wait for 100 ns; 
     
-------------------------------------------------------------------------
-- x80000000 < xFFFFFFF1
-- Expected value F= x00000001, CryOut= 0, Zero= 0,  overFlow =0
-------------------------------------------------------------------------
    s_A <= x"80000000";
    s_B <= x"FFFFFFF1";
    s_Opcode <= "110";
    wait for 100 ns; 

-------------------------------------------------------------------------
-- End of SLT test !!!!!
--  
--
-- 
--
--
--End of SLT Test !!!!!!
------------------------------------------------------------------------- 

-------------------------------------------------------------------------
-- Sub test !!!!!
--  
--
-- This will test our subfunction of our 32 bit ALU
--
--
--Sub Test
-------------------------------------------------------------------------

-------------------------------------------------------------------------
-- 0-0
-- Expected value F= x00000000, CryOut= 0, Zero= 1,  overFlow =0
-------------------------------------------------------------------------
    s_A <= x"00000000";
    s_B <= x"00000000";
    s_Opcode <= "111";
    wait for 100 ns;

-------------------------------------------------------------------------
-- 1-0
-- Expected value F= x00000001, CryOut= 0, Zero= 0,  overFlow =0
-------------------------------------------------------------------------
    s_A <= x"00000001";
    s_B <= x"00000000";
    s_Opcode <= "111";
    wait for 100 ns;

-------------------------------------------------------------------------
-- 0-1
-- Expected value F= xFFFFFFFF, CryOut= 0, Zero= 0,  overFlow =0
-------------------------------------------------------------------------
    s_A <= x"00000000";
    s_B <= x"00000001";
    s_Opcode <= "111";
    wait for 100 ns;

-------------------------------------------------------------------------
-- (-1)-(-1)
-- Expected value F= x00000000, CryOut= 0, Zero= 1,  overFlow =0
-------------------------------------------------------------------------
    s_A <= x"FFFFFFFF";
    s_B <= x"FFFFFFFF";
    s_Opcode <= "111";
    wait for 100 ns;

-------------------------------------------------------------------------
-- (-1)-(1)
-- Expected value F= xFFFFFFFD, CryOut= 0, Zero= 0,  overFlow =0
-------------------------------------------------------------------------
    s_A <= x"FFFFFFFF";
    s_B <= x"00000001";
    s_Opcode <= "111";
    wait for 100 ns;
     
-------------------------------------------------------------------------
-- 7FFFFFFF-(-2)
-- Expected value F= x80000002, CryOut= 0, Zero=0 ,  overFlow = 1
-------------------------------------------------------------------------
    s_A <= x"7FFFFFFF";
    s_B <= x"FFFFFFFD";
    s_Opcode <= "111";
    wait for 100 ns;

-------------------------------------------------------------------------
-- End of SUB test !!!!!
--  
--
-- 
--
--
--End of SUB Test !!!!!!
------------------------------------------------------------------------- 






  end process;
  
end behavioral;
