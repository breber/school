-------------------------------------------------------------------------
-- Group 9  :  Scott Connell, Brian Reber, Arjay Vander Velden
-- Project Part B
-- Due: November 9th, 2011
-------------------------------------------------------------------------

-- tb_control.vhd
-------------------------------------------------------------------------
-- DESCRIPTION:  This is the Control Logic testbench.
--               See the "Omniscient Spreadsheet" for more information
--               about what each instruction requires.
--               
-------------------------------------------------------------------------


library IEEE;
use IEEE.std_logic_1164.all;
use WORK.mips_package.all;


entity tb_control is

end tb_control;

architecture behavioral of tb_control is




Component Control_Logic is
  port(   instruction     :     in  std_logic_vector( 31 downto 0 );
          ALU_op          :     out std_logic_vector( 2 downto 0 );
          ALU_src         :     out std_logic;
          log_arith       :     out std_logic;
          leftOrRight     :     out std_logic;
          IsJump          :     out std_logic;
          IsBranch        :     out std_logic;
          RegWrite        :     out std_logic;
          MemWrite        :     out std_logic;
          MemRead         :     out std_logic;
          MemToReg        :     out std_logic_vector( 1 downto 0 );
          RegDest         :     out std_logic_vector( 1 downto 0 );
          W_H_B           :     out std_logic_vector( 2 downto 0 );
          WhichJB         :     out std_logic_vector( 3 downto 0 );
          shftAmount      :     out std_logic_vector( 1 downto 0 );
          isLui           :     out std_logic;
          NeedsLink       :     out std_logic   );
end component;
        



signal s_instruction                    : std_logic_vector( 31 downto 0 );
signal s_RegDest, s_MemToReg, s_shftAmount     : std_logic_vector( 1 downto 0 );
signal s_W_H_B, s_ALU_op     : std_logic_vector( 2 downto 0 );
signal s_ALU_src, s_log_arith, s_leftOrRight, s_IsJump, s_IsBranch, 
s_RegWrite, s_MemWrite ,s_MemRead, s_NeedsLink, s_isLui      : std_logic;   
signal s_WhichJB  : std_logic_vector( 3 downto 0 );                

begin
  testme: Control_Logic 

  port map(  instruction  => s_instruction,
             ALU_op       => s_ALU_op,
             ALU_src      => s_ALU_src,
             log_arith    => s_log_arith,
             leftOrRight  => s_leftOrRight,
             IsJump       => s_IsJump,
             IsBranch     => s_IsBranch,
             RegWrite     => s_RegWrite,
             MemWrite     => s_MemWrite,
             MemRead      => s_MemRead,
             MemToReg     => s_MemToReg,
             RegDest      => s_RegDest,
             W_H_B        => s_W_H_B,
             WhichJB      => s_WhichJB,
             shftAmount   => s_shftAmount,
             isLui        => s_isLui,
             NeedsLink    => s_NeedsLink);
  	        
  
process
begin


-------------------------------------------------------------------------
--add
-------------------------------------------------------------------------

s_instruction <= x"00000020";
wait for 100 ns;

-------------------------------------------------------------------------
--addi
-------------------------------------------------------------------------

s_instruction <= x"20000000";
wait for 100 ns;

-------------------------------------------------------------------------
--addiu
-------------------------------------------------------------------------

s_instruction <= x"24000000";
wait for 100 ns;

-------------------------------------------------------------------------
--addu
-------------------------------------------------------------------------

s_instruction <= x"00000021";
wait for 100 ns;

-------------------------------------------------------------------------
--and
-------------------------------------------------------------------------

s_instruction <= x"00000024";
wait for 100 ns;

-------------------------------------------------------------------------
--andi
-------------------------------------------------------------------------

s_instruction <= x"30000000";
wait for 100 ns;

-------------------------------------------------------------------------
--beq
-------------------------------------------------------------------------

s_instruction <= x"10000000";
wait for 100 ns;

-------------------------------------------------------------------------
--bgez
-------------------------------------------------------------------------

s_instruction <= x"04010000";
wait for 100 ns;

-------------------------------------------------------------------------
--bgezal
-------------------------------------------------------------------------

s_instruction <= x"04110000";
wait for 100 ns;

-------------------------------------------------------------------------
--bgtz
-------------------------------------------------------------------------

s_instruction <= x"1c000000";
wait for 100 ns;

-------------------------------------------------------------------------
--blez
-------------------------------------------------------------------------

s_instruction <= x"18000000";
wait for 100 ns;

-------------------------------------------------------------------------
--bltz
-------------------------------------------------------------------------

s_instruction <= x"04000000";
wait for 100 ns;

-------------------------------------------------------------------------
--bltzal
-------------------------------------------------------------------------

s_instruction <= x"04100000";
wait for 100 ns;

-------------------------------------------------------------------------
--bne
-------------------------------------------------------------------------

s_instruction <= x"14000000";
wait for 100 ns;

-------------------------------------------------------------------------
--j
-------------------------------------------------------------------------

s_instruction <= x"08000000";
wait for 100 ns;

-------------------------------------------------------------------------
--jal
-------------------------------------------------------------------------

s_instruction <= x"0c000000";
wait for 100 ns;

-------------------------------------------------------------------------
--jalr
-------------------------------------------------------------------------

s_instruction <= x"00000009";
wait for 100 ns;

-------------------------------------------------------------------------
--jr
-------------------------------------------------------------------------

s_instruction <= x"00000008";
wait for 100 ns;

-------------------------------------------------------------------------
--lb
-------------------------------------------------------------------------

s_instruction <= x"80000000";
wait for 100 ns;

-------------------------------------------------------------------------
--lbu
-------------------------------------------------------------------------

s_instruction <= x"90000000";
wait for 100 ns;

-------------------------------------------------------------------------
--lh
-------------------------------------------------------------------------

s_instruction <= x"84000000";
wait for 100 ns;

-------------------------------------------------------------------------
--lhu
-------------------------------------------------------------------------

s_instruction <= x"94000000";
wait for 100 ns;

-------------------------------------------------------------------------
--lui
-------------------------------------------------------------------------

s_instruction <= x"3c000000";
wait for 100 ns;

-------------------------------------------------------------------------
--lw
-------------------------------------------------------------------------

s_instruction <= x"8c000000";
wait for 100 ns;

-------------------------------------------------------------------------
--mul
-------------------------------------------------------------------------

s_instruction <= x"70000002";
wait for 100 ns;

-------------------------------------------------------------------------
--nor
-------------------------------------------------------------------------

s_instruction <= x"00000027";
wait for 100 ns;

-------------------------------------------------------------------------
--or
-------------------------------------------------------------------------

s_instruction <= x"00000025";
wait for 100 ns;

-------------------------------------------------------------------------
--ori
-------------------------------------------------------------------------

s_instruction <= x"34000000";
wait for 100 ns;

-------------------------------------------------------------------------
--sb
-------------------------------------------------------------------------

s_instruction <= x"a0000000";
wait for 100 ns;

-------------------------------------------------------------------------
--sh
-------------------------------------------------------------------------

s_instruction <= x"a4000000";
wait for 100 ns;


-------------------------------------------------------------------------
--sll
-------------------------------------------------------------------------

s_instruction <= x"00000000";
wait for 100 ns;

-------------------------------------------------------------------------
--sllv
-------------------------------------------------------------------------

s_instruction <= x"00000004";
wait for 100 ns;

-------------------------------------------------------------------------
--slt
-------------------------------------------------------------------------

s_instruction <= x"0000002a";
wait for 100 ns;

-------------------------------------------------------------------------
--slti
-------------------------------------------------------------------------

s_instruction <= x"28000000";
wait for 100 ns;

-------------------------------------------------------------------------
--sltiu
-------------------------------------------------------------------------

s_instruction <= x"2c000000";
wait for 100 ns;

-------------------------------------------------------------------------
--sltu
-------------------------------------------------------------------------

s_instruction <= x"0000002b";
wait for 100 ns;

-------------------------------------------------------------------------
--sra
-------------------------------------------------------------------------

s_instruction <= x"00000003";
wait for 100 ns;

-------------------------------------------------------------------------
--srav
-------------------------------------------------------------------------

s_instruction <= x"00000007";
wait for 100 ns;

-------------------------------------------------------------------------
--srl
-------------------------------------------------------------------------

s_instruction <= x"00000002";
wait for 100 ns;

-------------------------------------------------------------------------
--srlv
-------------------------------------------------------------------------

s_instruction <= x"00000006";
wait for 100 ns;

-------------------------------------------------------------------------
--sub
-------------------------------------------------------------------------

s_instruction <= x"00000022";
wait for 100 ns;

-------------------------------------------------------------------------
--subu
-------------------------------------------------------------------------

s_instruction <= x"00000023";
wait for 100 ns;

-------------------------------------------------------------------------
--sw
-------------------------------------------------------------------------

s_instruction <= x"ac000000";
wait for 100 ns;

-------------------------------------------------------------------------
--xor
-------------------------------------------------------------------------

s_instruction <= x"00000026";
wait for 100 ns;

-------------------------------------------------------------------------
--xori
-------------------------------------------------------------------------

s_instruction <= x"38000000";
wait for 100 ns;



end process;
  
end behavioral;




